`ifndef INSTMEM_V
`define INSTMEM_V

module INSTMEM(
    input[31:0] Addr,
    output[31:0] Inst
);
    wire[31:0] Rom[31:0];
    assign Rom[0]=32'b000000-00010-00011-00001-00000-100000;//add $1,$2,$3   $1=$2 + $3  
    assign Rom[1]=32'b000000-00010-00011-00001-00000-100010;//sub $1,$2,$3   $1=$2 - $3 
    assign Rom[2]=32'b000000-00010-00011-00001-00000-100100;//and $1,$2,$3   $1=$2 & $3
    assign Rom[3]=32'b000000-00010-00011-00001-00000-100101;//or $1,$2,$3    $1=$2 | $3 
    assign Rom[4]=32'b001000-00010-00001-0000000000001000;//addi $1,$2,1000 $1=$2+1000
	assign Rom[5]=32'b001100-00010-00001-0000000000001000;//andi $1,$2,1000  $1=$2 & 1000
    assign Rom[6]=32'b001101-00010-00001-0000000000001000;//ori $1,$2,1000   $1=$2 | 1000
    assign Rom[7]=32'b001111-00000-00001-0000000000000100;//lui $1,100     $1=100<<16//还未实现
    assign Rom[8]=32'b100011-00010-00001-0000000000000100;//lw $1,100($2)   $1=memory[$2 +10]
    assign Rom[9]=32'b101011-00010-00001-0000000000000100;//sw $1,100($2)    memory[$2+100]=$1 
    assign Rom[10]=32'b000100-00010-00001-0000000000000010;//beq $1,$2,10   if(Z==0) go to PC+4+10<<2
    assign Rom[11]=32'b000100-00010-00001-0000000000000010;//beq $1,$2,10   if(Z==1) dont go
    assign Rom[12]=32'b000101-00010-00001-0000000000000010;//bne $1,$2,10   if(Z==1) goto
    assign Rom[13]=32'b000101-00010-00001-0000000000000010;//bne $1,$2,10   if(Z==0) dont go
    assign Rom[14]=32'b000010-00000000000000000000010000;//j 10000        goto 10000

    assign Inst=Rom[Addr[6:2]];
endmodule
`endif