module DEC5T32E(I,En,Y);
    input[4:0] I;
    input En;
    output[31:0] Y;

	function[31:0] dec;
		input[4:0] I;
		input En;

		if(En)  
		    begin
		    case(I)
		    5'b0_0000 : dec = 32'b0000_0000_0000_0000_0000_0000_0000_0001 ;
		    5'b0_0001 : dec = 32'b0000_0000_0000_0000_0000_0000_0000_0010 ;
		    5'b0_0010 : dec = 32'b0000_0000_0000_0000_0000_0000_0000_0100 ;
			5'b0_0011 : dec = 32'b0000_0000_0000_0000_0000_0000_0000_1000 ;
			5'b0_0100 : dec = 32'b0000_0000_0000_0000_0000_0000_0001_0000 ;
			5'b0_0101 : dec = 32'b0000_0000_0000_0000_0000_0000_0010_0000 ;
			5'b0_0110 : dec = 32'b0000_0000_0000_0000_0000_0000_0100_0000 ;
			5'b0_0111 : dec = 32'b0000_0000_0000_0000_0000_0000_1000_0000 ;
			5'b0_1000 : dec = 32'b0000_0000_0000_0000_0000_0001_0000_0000 ;
			5'b0_1001 : dec = 32'b0000_0000_0000_0000_0000_0010_0000_0000 ;
			5'b0_1010 : dec = 32'b0000_0000_0000_0000_0000_0100_0000_0000 ;
			5'b0_1011 : dec = 32'b0000_0000_0000_0000_0000_1000_0000_0000 ;
			5'b0_1100 : dec = 32'b0000_0000_0000_0000_0001_0000_0000_0000 ;
			5'b0_1101 : dec = 32'b0000_0000_0000_0000_0010_0000_0000_0000 ;
			5'b0_1110 : dec = 32'b0000_0000_0000_0000_0100_0000_0000_0000 ;
			5'b0_1111 : dec = 32'b0000_0000_0000_0000_1000_0000_0000_0000 ;
			5'b1_0000 : dec = 32'b0000_0000_0000_0001_0000_0000_0000_0000 ;
			5'b1_0001 : dec = 32'b0000_0000_0000_0010_0000_0000_0000_0000 ;
			5'b1_0010 : dec = 32'b0000_0000_0000_0100_0000_0000_0000_0000 ;
			5'b1_0011 : dec = 32'b0000_0000_0000_1000_0000_0000_0000_0000 ;
			5'b1_0100 : dec = 32'b0000_0000_0001_0000_0000_0000_0000_0000 ;
			5'b1_0101 : dec = 32'b0000_0000_0010_0000_0000_0000_0000_0000 ;
			5'b1_0110 : dec = 32'b0000_0000_0100_0000_0000_0000_0000_0000 ;
			5'b1_0111 : dec = 32'b0000_0000_1000_0000_0000_0000_0000_0000 ;
			5'b1_1000 : dec = 32'b0000_0001_0000_0000_0000_0000_0000_0000 ;
		    5'b1_1001 : dec = 32'b0000_0010_0000_0000_0000_0000_0000_0000 ;
			5'b1_1010 : dec = 32'b0000_0100_0000_0000_0000_0000_0000_0000 ;
			5'b1_1011 : dec = 32'b0000_1000_0000_0000_0000_0000_0000_0000 ;
			5'b1_1100 : dec = 32'b0001_0000_0000_0000_0000_0000_0000_0000 ;
			5'b1_1101 : dec = 32'b0010_0000_0000_0000_0000_0000_0000_0000 ;
		    5'b1_1110 : dec = 32'b0100_0000_0000_0000_0000_0000_0000_0000 ;
			5'b1_1111 : dec = 32'b1000_0000_0000_0000_0000_0000_0000_0000 ;
			default   : dec = 32'b0000_0000_0000_0000_0000_0000_0000_0000 ;
            endcase
		    end
    	else  dec = 32'b0000_0000_0000_0000_0000_0000_0000_0000 ;
	endfunction

	assign Y=dec(I,En);
endmodule